-- Copyright (C) 2022  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and any partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details, at
-- https://fpgasoftware.intel.com/eula.

-- PROGRAM		"Quartus Prime"
-- VERSION		"Version 21.1.1 Build 850 06/23/2022 SJ Lite Edition"
-- CREATED		"Wed Nov  5 20:45:45 2025"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY BCD_COUNTER IS 
	PORT
	(
		clk :  IN  STD_LOGIC;
		CLRN :  IN  STD_LOGIC;
		Q0 :  OUT  STD_LOGIC;
		Q1 :  OUT  STD_LOGIC;
		Q2 :  OUT  STD_LOGIC;
		Q3 :  OUT  STD_LOGIC
	);
END BCD_COUNTER;

ARCHITECTURE bdf_type OF BCD_COUNTER IS 

SIGNAL	SYNTHESIZED_WIRE_22 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_1 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_2 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_3 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_23 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_24 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_4 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_25 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_7 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_8 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_9 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_26 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_27 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_12 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_13 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_14 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_15 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_16 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_17 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_18 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_19 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_21 :  STD_LOGIC;


BEGIN 
Q0 <= SYNTHESIZED_WIRE_23;
Q1 <= SYNTHESIZED_WIRE_24;
Q2 <= SYNTHESIZED_WIRE_25;
Q3 <= SYNTHESIZED_WIRE_27;
SYNTHESIZED_WIRE_1 <= '1';
SYNTHESIZED_WIRE_3 <= '1';
SYNTHESIZED_WIRE_15 <= '1';
SYNTHESIZED_WIRE_17 <= '1';



PROCESS(CLRN,clk,SYNTHESIZED_WIRE_1)
BEGIN
IF (clk = '0') THEN
	SYNTHESIZED_WIRE_23 <= '0';
ELSIF (SYNTHESIZED_WIRE_1 = '0') THEN
	SYNTHESIZED_WIRE_23 <= '1';
ELSIF (RISING_EDGE(CLRN)) THEN
	SYNTHESIZED_WIRE_23 <= SYNTHESIZED_WIRE_22;
END IF;
END PROCESS;


PROCESS(CLRN,clk,SYNTHESIZED_WIRE_3)
BEGIN
IF (clk = '0') THEN
	SYNTHESIZED_WIRE_24 <= '0';
ELSIF (SYNTHESIZED_WIRE_3 = '0') THEN
	SYNTHESIZED_WIRE_24 <= '1';
ELSIF (RISING_EDGE(CLRN)) THEN
	SYNTHESIZED_WIRE_24 <= SYNTHESIZED_WIRE_2;
END IF;
END PROCESS;


SYNTHESIZED_WIRE_9 <= SYNTHESIZED_WIRE_23 AND SYNTHESIZED_WIRE_24 AND SYNTHESIZED_WIRE_4;


SYNTHESIZED_WIRE_12 <= SYNTHESIZED_WIRE_23 AND SYNTHESIZED_WIRE_24 AND SYNTHESIZED_WIRE_25;


SYNTHESIZED_WIRE_18 <= SYNTHESIZED_WIRE_22 AND SYNTHESIZED_WIRE_24;


SYNTHESIZED_WIRE_7 <= SYNTHESIZED_WIRE_22 AND SYNTHESIZED_WIRE_25;


SYNTHESIZED_WIRE_14 <= SYNTHESIZED_WIRE_7 OR SYNTHESIZED_WIRE_8 OR SYNTHESIZED_WIRE_9;


SYNTHESIZED_WIRE_8 <= SYNTHESIZED_WIRE_26 AND SYNTHESIZED_WIRE_25;


SYNTHESIZED_WIRE_13 <= SYNTHESIZED_WIRE_22 AND SYNTHESIZED_WIRE_27;


SYNTHESIZED_WIRE_16 <= SYNTHESIZED_WIRE_12 OR SYNTHESIZED_WIRE_13;



PROCESS(CLRN,clk,SYNTHESIZED_WIRE_15)
BEGIN
IF (clk = '0') THEN
	SYNTHESIZED_WIRE_25 <= '0';
ELSIF (SYNTHESIZED_WIRE_15 = '0') THEN
	SYNTHESIZED_WIRE_25 <= '1';
ELSIF (RISING_EDGE(CLRN)) THEN
	SYNTHESIZED_WIRE_25 <= SYNTHESIZED_WIRE_14;
END IF;
END PROCESS;





PROCESS(CLRN,clk,SYNTHESIZED_WIRE_17)
BEGIN
IF (clk = '0') THEN
	SYNTHESIZED_WIRE_27 <= '0';
ELSIF (SYNTHESIZED_WIRE_17 = '0') THEN
	SYNTHESIZED_WIRE_27 <= '1';
ELSIF (RISING_EDGE(CLRN)) THEN
	SYNTHESIZED_WIRE_27 <= SYNTHESIZED_WIRE_16;
END IF;
END PROCESS;


SYNTHESIZED_WIRE_22 <= NOT(SYNTHESIZED_WIRE_23);



SYNTHESIZED_WIRE_26 <= NOT(SYNTHESIZED_WIRE_24);



SYNTHESIZED_WIRE_4 <= NOT(SYNTHESIZED_WIRE_25);



SYNTHESIZED_WIRE_21 <= NOT(SYNTHESIZED_WIRE_27);



SYNTHESIZED_WIRE_2 <= SYNTHESIZED_WIRE_18 OR SYNTHESIZED_WIRE_19;


SYNTHESIZED_WIRE_19 <= SYNTHESIZED_WIRE_23 AND SYNTHESIZED_WIRE_26 AND SYNTHESIZED_WIRE_21;


END bdf_type;